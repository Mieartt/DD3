library ieee;
use ieee.std_logic_116.all;
entity abdou is
port ( wednin, khcham   : in std_logic;
        fom             : out std_logic);
end entity;
architecture behavior of abdou is
signal sch3ar   : std_logic_vector (2 downto 0);
signal jel : std_logic;
begin
ch3ar <= jel;
end architecture;