library ieee;
use ieee.std_logic_116.all;
entity abdou is
port ( wednin, khcham : in std_logic;
        fom           : out std_logic);
end entity;